library verilog;
use verilog.vl_types.all;
entity upc_check_testbench is
end upc_check_testbench;
