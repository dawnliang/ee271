library verilog;
use verilog.vl_types.all;
entity upc_check_display_testbench is
end upc_check_display_testbench;
