library verilog;
use verilog.vl_types.all;
entity upc_display_testbench is
end upc_display_testbench;
